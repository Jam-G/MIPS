library verilog;
use verilog.vl_types.all;
entity ID_EX is
    port(
        Clk             : in     vl_logic;
        stall           : in     vl_logic;
        flush           : in     vl_logic;
        PC_4_ID         : in     vl_logic_vector(31 downto 0);
        op_ID           : in     vl_logic_vector(5 downto 0);
        Condition_ID    : in     vl_logic_vector(2 downto 0);
        Branch_ID       : in     vl_logic;
        MemWrite_ID     : in     vl_logic;
        RegWrite_ID     : in     vl_logic;
        MemRead_ID      : in     vl_logic;
        Jump_ID         : in     vl_logic;
        ExResultSrc_ID  : in     vl_logic_vector(1 downto 0);
        ALUSrcA_ID      : in     vl_logic;
        ALUSrcB_ID      : in     vl_logic;
        ALUop_ID        : in     vl_logic_vector(3 downto 0);
        regdst_ID       : in     vl_logic_vector(1 downto 0);
        ShiftAmountSrc_ID: in     vl_logic;
        ShiftOp_ID      : in     vl_logic_vector(1 downto 0);
        A_in_ID         : in     vl_logic_vector(31 downto 0);
        B_in_ID         : in     vl_logic_vector(31 downto 0);
        Rs_ID           : in     vl_logic_vector(4 downto 0);
        Rt_ID           : in     vl_logic_vector(4 downto 0);
        Rd_ID           : in     vl_logic_vector(4 downto 0);
        Immediate32_ID  : in     vl_logic_vector(31 downto 0);
        Shamt_ID        : in     vl_logic_vector(4 downto 0);
        loaduse_in      : in     vl_logic;
        PC_4_EX         : out    vl_logic_vector(31 downto 0);
        op_EX           : out    vl_logic_vector(5 downto 0);
        Condition_EX    : out    vl_logic_vector(2 downto 0);
        Branch_EX       : out    vl_logic;
        MemWrite_EX     : out    vl_logic;
        RegWrite_EX     : out    vl_logic;
        MemRead_EX      : out    vl_logic;
        Jump_EX         : out    vl_logic;
        ExResultSrc_EX  : out    vl_logic_vector(1 downto 0);
        ALUSrcA_EX      : out    vl_logic;
        ALUSrcB_EX      : out    vl_logic;
        ALUop_EX        : out    vl_logic_vector(3 downto 0);
        regdst_EX       : out    vl_logic_vector(1 downto 0);
        ShiftAmountSrc_EX: out    vl_logic;
        ShiftOp_EX      : out    vl_logic_vector(1 downto 0);
        A_in_EX         : out    vl_logic_vector(31 downto 0);
        B_in_EX         : out    vl_logic_vector(31 downto 0);
        Rs_EX           : out    vl_logic_vector(4 downto 0);
        Rt_EX           : out    vl_logic_vector(4 downto 0);
        Rd_EX           : out    vl_logic_vector(4 downto 0);
        Immediate32_EX  : out    vl_logic_vector(31 downto 0);
        Shamt_EX        : out    vl_logic_vector(4 downto 0);
        loaduse_out     : out    vl_logic
    );
end ID_EX;
