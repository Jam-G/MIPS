library verilog;
use verilog.vl_types.all;
entity Pipeline_vlg_tst is
end Pipeline_vlg_tst;
